_.vhdl