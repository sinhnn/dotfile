--------------------------------------------------------------------------------
-- Project name   :
-- File name      : !!FILE
-- Created date   : !!DATE
-- Author         : Ngoc-Sinh Nguyen
-- Last modified  : !!DATE
-- Desc           :
--------------------------------------------------------------------------------

